LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.ALL;

PACKAGE parameter IS
  CONSTANT SIGNAL_WIDTH :INTEGER := 16;
  --CONSTANT REGISTER_LENGTH : INTEGER := 10000;
  CONSTANT xcorr_SIGNAL_WIDTH : INTEGER := 32;
  CONSTANT xcorr_MAXLAG : INTEGER := 140;
  CONSTANT LEN_DATA: integer:=23;
  CONSTANT POWER_WINDOW : INTEGER := 100;
  CONSTANT xcorr_WINDOW : INTEGER := 10000;
  
  TYPE outputdata IS ARRAY (0 TO 1) OF STD_LOGIC_VECTOR(SIGNAL_WIDTH-1 DOWNTO 0);
  TYPE xcorrdata IS ARRAY (0 TO 2*xcorr_MAXLAG-1) OF STD_LOGIC_VECTOR(xcorr_SIGNAL_WIDTH-1 DOWNTO 0);
  
  
END PACKAGE;

